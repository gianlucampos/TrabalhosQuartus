--**************************************--
--			Morgana M.A.R.
--**************************************--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

ENTITY Raiz IS
	PORT(
			CLOCK_50: IN STD_LOGIC;
			SW		: IN STD_LOGIC_VECTOR (7 downto 0 ); --Interruptores 
			BUTTON	: IN STD_LOGIC_VECTOR (2 downto 0 ); --Botao 3
			HEX3_D	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX2_D	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX1_D	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX0_D	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
			);END Raiz;

ARCHITECTURE comportamento OF Raiz IS
SIGNAL OUT_Raiz			: STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL saida_display	: STD_LOGIC_VECTOR (15 downto 0);
begin
process(CLOCK_50)
	variable r: std_logic_vector(3 downto 0);
	variable d: std_logic_vector(4 downto 0);
	variable s, temp: std_logic_vector(8 downto 0);
	begin
		if CLOCK_50'event and CLOCK_50 = '1' then
				if BUTTON(0) ='0' then
					r:="0001";
					d:="00010";
					s:="000000100";
				else 
					temp := SW(7 downto 0)-s;
					if (temp(8)='0')then
						r:=r+1;
						d:=d+2;
						s:=s+d+1;
					else 
						OUT_Raiz <= "000000000000"&r;
					end if;
				end if;				
		end if;
end process;
PROCESS (CLOCK_50)
BEGIN
	IF CLOCK_50'event and CLOCK_50='1'  THEN
	saida_display <= OUT_Raiz(15 DOWNTO 0);
CASE saida_display IS
WHEN "0000000000000000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--0
WHEN "0000000000000001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--1
WHEN "0000000000000010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--2
WHEN "0000000000000011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--3
WHEN "0000000000000100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--4
WHEN "0000000000000101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--5
WHEN "0000000000000110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--6
WHEN "0000000000000111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--7
WHEN "0000000000001000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--8
WHEN "0000000000001001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--9
WHEN "0000000000001010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--10
WHEN "0000000000001011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--11
WHEN "0000000000001100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--12
WHEN "0000000000001101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--13
WHEN "0000000000001110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--14
WHEN "0000000000001111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--15
WHEN "0000000000010000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--16
WHEN "0000000000010001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--17
WHEN "0000000000010010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--18
WHEN "0000000000010011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--19
WHEN "0000000000010100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--20
WHEN "0000000000010101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--21
WHEN "0000000000010110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--22
WHEN "0000000000010111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--23
WHEN "0000000000011000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--24
WHEN "0000000000011001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--25
WHEN "0000000000011010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--26
WHEN "0000000000011011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--27
WHEN "0000000000011100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--28
WHEN "0000000000011101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--29
WHEN "0000000000011110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--30
WHEN "0000000000011111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--31
WHEN "0000000000100000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--32
WHEN "0000000000100001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--33
WHEN "0000000000100010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--34
WHEN "0000000000100011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--35
WHEN "0000000000100100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--36
WHEN "0000000000100101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--37
WHEN "0000000000100110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--38
WHEN "0000000000100111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--39
WHEN "0000000000101000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--40
WHEN "0000000000101001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--41
WHEN "0000000000101010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--42
WHEN "0000000000101011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--43
WHEN "0000000000101100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--44
WHEN "0000000000101101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--45
WHEN "0000000000101110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--46
WHEN "0000000000101111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--47
WHEN "0000000000110000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--48
WHEN "0000000000110001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--49
WHEN "0000000000110010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--50
WHEN "0000000000110011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--51
WHEN "0000000000110100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--52
WHEN "0000000000110101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--53
WHEN "0000000000110110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--54
WHEN "0000000000110111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--55
WHEN "0000000000111000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--56
WHEN "0000000000111001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--57
WHEN "0000000000111010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--58
WHEN "0000000000111011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--59
WHEN "0000000000111100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--60
WHEN "0000000000111101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--61
WHEN "0000000000111110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--62
WHEN "0000000000111111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--63
WHEN "0000000001000000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--64
WHEN "0000000001000001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--65
WHEN "0000000001000010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--66
WHEN "0000000001000011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--67
WHEN "0000000001000100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--68
WHEN "0000000001000101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--69
WHEN "0000000001000110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--70
WHEN "0000000001000111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--71
WHEN "0000000001001000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--72
WHEN "0000000001001001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--73
WHEN "0000000001001010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--74
WHEN "0000000001001011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--75
WHEN "0000000001001100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--76
WHEN "0000000001001101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--77
WHEN "0000000001001110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--78
WHEN "0000000001001111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--79
WHEN "0000000001010000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--80
WHEN "0000000001010001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--81
WHEN "0000000001010010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--82
WHEN "0000000001010011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--83
WHEN "0000000001010100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--84
WHEN "0000000001010101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--85
WHEN "0000000001010110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--86
WHEN "0000000001010111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--87
WHEN "0000000001011000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--88
WHEN "0000000001011001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--89
WHEN "0000000001011010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--90
WHEN "0000000001011011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--91
WHEN "0000000001011100" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--92
WHEN "0000000001011101" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--93
WHEN "0000000001011110" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--94
WHEN "0000000001011111" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--95
WHEN "0000000001100000" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--96
WHEN "0000000001100001" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--97
WHEN "0000000001100010" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--98
WHEN "0000000001100011" => HEX3_D <= "1000000"; HEX2_D <= "1000000"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--99
WHEN "0000000001100100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--100
WHEN "0000000001100101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--101
WHEN "0000000001100110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--102
WHEN "0000000001100111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--103
WHEN "0000000001101000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--104
WHEN "0000000001101001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--105
WHEN "0000000001101010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--106
WHEN "0000000001101011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--107
WHEN "0000000001101100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--108
WHEN "0000000001101101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--109
WHEN "0000000001101110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--110
WHEN "0000000001101111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--111
WHEN "0000000001110000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--112
WHEN "0000000001110001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--113
WHEN "0000000001110010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--114
WHEN "0000000001110011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--115
WHEN "0000000001110100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--116
WHEN "0000000001110101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--117
WHEN "0000000001110110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--118
WHEN "0000000001110111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--119
WHEN "0000000001111000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--120
WHEN "0000000001111001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--121
WHEN "0000000001111010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--122
WHEN "0000000001111011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--123
WHEN "0000000001111100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--124
WHEN "0000000001111101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--125
WHEN "0000000001111110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--126
WHEN "0000000001111111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--127
WHEN "0000000010000000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--128
WHEN "0000000010000001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--129
WHEN "0000000010000010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--130
WHEN "0000000010000011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--131
WHEN "0000000010000100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--132
WHEN "0000000010000101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--133
WHEN "0000000010000110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--134
WHEN "0000000010000111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--135
WHEN "0000000010001000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--136
WHEN "0000000010001001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--137
WHEN "0000000010001010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--138
WHEN "0000000010001011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--139
WHEN "0000000010001100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--140
WHEN "0000000010001101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--141
WHEN "0000000010001110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--142
WHEN "0000000010001111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--143
WHEN "0000000010010000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--144
WHEN "0000000010010001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--145
WHEN "0000000010010010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--146
WHEN "0000000010010011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--147
WHEN "0000000010010100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--148
WHEN "0000000010010101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--149
WHEN "0000000010010110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--150
WHEN "0000000010010111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--151
WHEN "0000000010011000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--152
WHEN "0000000010011001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--153
WHEN "0000000010011010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--154
WHEN "0000000010011011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--155
WHEN "0000000010011100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--156
WHEN "0000000010011101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--157
WHEN "0000000010011110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--158
WHEN "0000000010011111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--159
WHEN "0000000010100000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--160
WHEN "0000000010100001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--161
WHEN "0000000010100010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--162
WHEN "0000000010100011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--163
WHEN "0000000010100100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--164
WHEN "0000000010100101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--165
WHEN "0000000010100110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--166
WHEN "0000000010100111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--167
WHEN "0000000010101000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--168
WHEN "0000000010101001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--169
WHEN "0000000010101010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--170
WHEN "0000000010101011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--171
WHEN "0000000010101100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--172
WHEN "0000000010101101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--173
WHEN "0000000010101110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--174
WHEN "0000000010101111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--175
WHEN "0000000010110000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--176
WHEN "0000000010110001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--177
WHEN "0000000010110010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--178
WHEN "0000000010110011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--179
WHEN "0000000010110100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--180
WHEN "0000000010110101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--181
WHEN "0000000010110110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--182
WHEN "0000000010110111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--183
WHEN "0000000010111000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--184
WHEN "0000000010111001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--185
WHEN "0000000010111010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--186
WHEN "0000000010111011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--187
WHEN "0000000010111100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--188
WHEN "0000000010111101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--189
WHEN "0000000010111110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--190
WHEN "0000000010111111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--191
WHEN "0000000011000000" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--192
WHEN "0000000011000001" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--193
WHEN "0000000011000010" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--194
WHEN "0000000011000011" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--195
WHEN "0000000011000100" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--196
WHEN "0000000011000101" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--197
WHEN "0000000011000110" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--198
WHEN "0000000011000111" => HEX3_D <= "1000000"; HEX2_D <= "1111001"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--199
WHEN "0000000011001000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--200
WHEN "0000000011001001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--201
WHEN "0000000011001010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--202
WHEN "0000000011001011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--203
WHEN "0000000011001100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--204
WHEN "0000000011001101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--205
WHEN "0000000011001110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--206
WHEN "0000000011001111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--207
WHEN "0000000011010000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--208
WHEN "0000000011010001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--209
WHEN "0000000011010010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--210
WHEN "0000000011010011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--211
WHEN "0000000011010100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--212
WHEN "0000000011010101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--213
WHEN "0000000011010110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--214
WHEN "0000000011010111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--215
WHEN "0000000011011000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--216
WHEN "0000000011011001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--217
WHEN "0000000011011010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--218
WHEN "0000000011011011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--219
WHEN "0000000011011100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--220
WHEN "0000000011011101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--221
WHEN "0000000011011110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--222
WHEN "0000000011011111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--223
WHEN "0000000011100000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--224
WHEN "0000000011100001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--225
WHEN "0000000011100010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--226
WHEN "0000000011100011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--227
WHEN "0000000011100100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--228
WHEN "0000000011100101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--229
WHEN "0000000011100110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--230
WHEN "0000000011100111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--231
WHEN "0000000011101000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--232
WHEN "0000000011101001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--233
WHEN "0000000011101010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--234
WHEN "0000000011101011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--235
WHEN "0000000011101100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--236
WHEN "0000000011101101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--237
WHEN "0000000011101110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--238
WHEN "0000000011101111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--239
WHEN "0000000011110000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--240
WHEN "0000000011110001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--241
WHEN "0000000011110010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--242
WHEN "0000000011110011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--243
WHEN "0000000011110100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--244
WHEN "0000000011110101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--245
WHEN "0000000011110110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--246
WHEN "0000000011110111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--247
WHEN "0000000011111000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--248
WHEN "0000000011111001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--249
WHEN "0000000011111010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--250
WHEN "0000000011111011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--251
WHEN "0000000011111100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--252
WHEN "0000000011111101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--253
WHEN "0000000011111110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--254
WHEN "0000000011111111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--255
WHEN "0000000100000000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--256
WHEN "0000000100000001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--257
WHEN "0000000100000010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--258
WHEN "0000000100000011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--259
WHEN "0000000100000100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--260
WHEN "0000000100000101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--261
WHEN "0000000100000110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--262
WHEN "0000000100000111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--263
WHEN "0000000100001000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--264
WHEN "0000000100001001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--265
WHEN "0000000100001010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--266
WHEN "0000000100001011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--267
WHEN "0000000100001100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--268
WHEN "0000000100001101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--269
WHEN "0000000100001110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--270
WHEN "0000000100001111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--271
WHEN "0000000100010000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--272
WHEN "0000000100010001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--273
WHEN "0000000100010010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--274
WHEN "0000000100010011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--275
WHEN "0000000100010100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--276
WHEN "0000000100010101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--277
WHEN "0000000100010110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--278
WHEN "0000000100010111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--279
WHEN "0000000100011000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--280
WHEN "0000000100011001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--281
WHEN "0000000100011010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--282
WHEN "0000000100011011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--283
WHEN "0000000100011100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--284
WHEN "0000000100011101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--285
WHEN "0000000100011110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--286
WHEN "0000000100011111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--287
WHEN "0000000100100000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--288
WHEN "0000000100100001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--289
WHEN "0000000100100010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--290
WHEN "0000000100100011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--291
WHEN "0000000100100100" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--292
WHEN "0000000100100101" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--293
WHEN "0000000100100110" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--294
WHEN "0000000100100111" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--295
WHEN "0000000100101000" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--296
WHEN "0000000100101001" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--297
WHEN "0000000100101010" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--298
WHEN "0000000100101011" => HEX3_D <= "1000000"; HEX2_D <= "0100100"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--299
WHEN "0000000100101100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--300
WHEN "0000000100101101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--301
WHEN "0000000100101110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--302
WHEN "0000000100101111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--303
WHEN "0000000100110000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--304
WHEN "0000000100110001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--305
WHEN "0000000100110010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--306
WHEN "0000000100110011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--307
WHEN "0000000100110100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--308
WHEN "0000000100110101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--309
WHEN "0000000100110110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--310
WHEN "0000000100110111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--311
WHEN "0000000100111000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--312
WHEN "0000000100111001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--313
WHEN "0000000100111010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--314
WHEN "0000000100111011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--315
WHEN "0000000100111100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--316
WHEN "0000000100111101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--317
WHEN "0000000100111110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--318
WHEN "0000000100111111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--319
WHEN "0000000101000000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--320
WHEN "0000000101000001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--321
WHEN "0000000101000010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--322
WHEN "0000000101000011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--323
WHEN "0000000101000100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--324
WHEN "0000000101000101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--325
WHEN "0000000101000110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--326
WHEN "0000000101000111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--327
WHEN "0000000101001000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--328
WHEN "0000000101001001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--329
WHEN "0000000101001010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--330
WHEN "0000000101001011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--331
WHEN "0000000101001100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--332
WHEN "0000000101001101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--333
WHEN "0000000101001110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--334
WHEN "0000000101001111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--335
WHEN "0000000101010000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--336
WHEN "0000000101010001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--337
WHEN "0000000101010010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--338
WHEN "0000000101010011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--339
WHEN "0000000101010100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--340
WHEN "0000000101010101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--341
WHEN "0000000101010110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--342
WHEN "0000000101010111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--343
WHEN "0000000101011000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--344
WHEN "0000000101011001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--345
WHEN "0000000101011010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--346
WHEN "0000000101011011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--347
WHEN "0000000101011100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--348
WHEN "0000000101011101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--349
WHEN "0000000101011110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--350
WHEN "0000000101011111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--351
WHEN "0000000101100000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--352
WHEN "0000000101100001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--353
WHEN "0000000101100010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--354
WHEN "0000000101100011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--355
WHEN "0000000101100100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--356
WHEN "0000000101100101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--357
WHEN "0000000101100110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--358
WHEN "0000000101100111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--359
WHEN "0000000101101000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--360
WHEN "0000000101101001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--361
WHEN "0000000101101010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--362
WHEN "0000000101101011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--363
WHEN "0000000101101100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--364
WHEN "0000000101101101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--365
WHEN "0000000101101110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--366
WHEN "0000000101101111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--367
WHEN "0000000101110000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--368
WHEN "0000000101110001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--369
WHEN "0000000101110010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--370
WHEN "0000000101110011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--371
WHEN "0000000101110100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--372
WHEN "0000000101110101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--373
WHEN "0000000101110110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--374
WHEN "0000000101110111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--375
WHEN "0000000101111000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--376
WHEN "0000000101111001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--377
WHEN "0000000101111010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--378
WHEN "0000000101111011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--379
WHEN "0000000101111100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--380
WHEN "0000000101111101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--381
WHEN "0000000101111110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--382
WHEN "0000000101111111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--383
WHEN "0000000110000000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--384
WHEN "0000000110000001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--385
WHEN "0000000110000010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--386
WHEN "0000000110000011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--387
WHEN "0000000110000100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--388
WHEN "0000000110000101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--389
WHEN "0000000110000110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--390
WHEN "0000000110000111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--391
WHEN "0000000110001000" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--392
WHEN "0000000110001001" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--393
WHEN "0000000110001010" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--394
WHEN "0000000110001011" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--395
WHEN "0000000110001100" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--396
WHEN "0000000110001101" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--397
WHEN "0000000110001110" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--398
WHEN "0000000110001111" => HEX3_D <= "1000000"; HEX2_D <= "0110000"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--399
WHEN "0000000110010000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--400
WHEN "0000000110010001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--401
WHEN "0000000110010010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--402
WHEN "0000000110010011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--403
WHEN "0000000110010100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--404
WHEN "0000000110010101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--405
WHEN "0000000110010110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--406
WHEN "0000000110010111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--407
WHEN "0000000110011000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--408
WHEN "0000000110011001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--409
WHEN "0000000110011010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--410
WHEN "0000000110011011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--411
WHEN "0000000110011100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--412
WHEN "0000000110011101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--413
WHEN "0000000110011110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--414
WHEN "0000000110011111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--415
WHEN "0000000110100000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--416
WHEN "0000000110100001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--417
WHEN "0000000110100010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--418
WHEN "0000000110100011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--419
WHEN "0000000110100100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--420
WHEN "0000000110100101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--421
WHEN "0000000110100110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--422
WHEN "0000000110100111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--423
WHEN "0000000110101000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--424
WHEN "0000000110101001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--425
WHEN "0000000110101010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--426
WHEN "0000000110101011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--427
WHEN "0000000110101100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--428
WHEN "0000000110101101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--429
WHEN "0000000110101110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--430
WHEN "0000000110101111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--431
WHEN "0000000110110000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--432
WHEN "0000000110110001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--433
WHEN "0000000110110010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--434
WHEN "0000000110110011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--435
WHEN "0000000110110100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--436
WHEN "0000000110110101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--437
WHEN "0000000110110110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--438
WHEN "0000000110110111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--439
WHEN "0000000110111000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--440
WHEN "0000000110111001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--441
WHEN "0000000110111010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--442
WHEN "0000000110111011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--443
WHEN "0000000110111100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--444
WHEN "0000000110111101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--445
WHEN "0000000110111110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--446
WHEN "0000000110111111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--447
WHEN "0000000111000000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--448
WHEN "0000000111000001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--449
WHEN "0000000111000010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--450
WHEN "0000000111000011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--451
WHEN "0000000111000100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--452
WHEN "0000000111000101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--453
WHEN "0000000111000110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--454
WHEN "0000000111000111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--455
WHEN "0000000111001000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--456
WHEN "0000000111001001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--457
WHEN "0000000111001010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--458
WHEN "0000000111001011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--459
WHEN "0000000111001100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--460
WHEN "0000000111001101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--461
WHEN "0000000111001110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--462
WHEN "0000000111001111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--463
WHEN "0000000111010000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--464
WHEN "0000000111010001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--465
WHEN "0000000111010010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--466
WHEN "0000000111010011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--467
WHEN "0000000111010100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--468
WHEN "0000000111010101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--469
WHEN "0000000111010110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--470
WHEN "0000000111010111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--471
WHEN "0000000111011000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--472
WHEN "0000000111011001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--473
WHEN "0000000111011010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--474
WHEN "0000000111011011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--475
WHEN "0000000111011100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--476
WHEN "0000000111011101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--477
WHEN "0000000111011110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--478
WHEN "0000000111011111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--479
WHEN "0000000111100000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--480
WHEN "0000000111100001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--481
WHEN "0000000111100010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--482
WHEN "0000000111100011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--483
WHEN "0000000111100100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--484
WHEN "0000000111100101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--485
WHEN "0000000111100110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--486
WHEN "0000000111100111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--487
WHEN "0000000111101000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--488
WHEN "0000000111101001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--489
WHEN "0000000111101010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--490
WHEN "0000000111101011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--491
WHEN "0000000111101100" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--492
WHEN "0000000111101101" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--493
WHEN "0000000111101110" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--494
WHEN "0000000111101111" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--495
WHEN "0000000111110000" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--496
WHEN "0000000111110001" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--497
WHEN "0000000111110010" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--498
WHEN "0000000111110011" => HEX3_D <= "1000000"; HEX2_D <= "0011001"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--499
WHEN "0000000111110100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--500
WHEN "0000000111110101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--501
WHEN "0000000111110110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--502
WHEN "0000000111110111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--503
WHEN "0000000111111000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--504
WHEN "0000000111111001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--505
WHEN "0000000111111010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--506
WHEN "0000000111111011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--507
WHEN "0000000111111100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--508
WHEN "0000000111111101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--509
WHEN "0000000111111110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--510
WHEN "0000000111111111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--511
WHEN "0000001000000000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--512
WHEN "0000001000000001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--513
WHEN "0000001000000010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--514
WHEN "0000001000000011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--515
WHEN "0000001000000100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--516
WHEN "0000001000000101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--517
WHEN "0000001000000110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--518
WHEN "0000001000000111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--519
WHEN "0000001000001000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--520
WHEN "0000001000001001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--521
WHEN "0000001000001010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--522
WHEN "0000001000001011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--523
WHEN "0000001000001100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--524
WHEN "0000001000001101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--525
WHEN "0000001000001110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--526
WHEN "0000001000001111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--527
WHEN "0000001000010000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--528
WHEN "0000001000010001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--529
WHEN "0000001000010010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--530
WHEN "0000001000010011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--531
WHEN "0000001000010100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--532
WHEN "0000001000010101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--533
WHEN "0000001000010110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--534
WHEN "0000001000010111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--535
WHEN "0000001000011000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--536
WHEN "0000001000011001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--537
WHEN "0000001000011010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--538
WHEN "0000001000011011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--539
WHEN "0000001000011100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--540
WHEN "0000001000011101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--541
WHEN "0000001000011110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--542
WHEN "0000001000011111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--543
WHEN "0000001000100000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--544
WHEN "0000001000100001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--545
WHEN "0000001000100010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--546
WHEN "0000001000100011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--547
WHEN "0000001000100100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--548
WHEN "0000001000100101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--549
WHEN "0000001000100110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--550
WHEN "0000001000100111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--551
WHEN "0000001000101000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--552
WHEN "0000001000101001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--553
WHEN "0000001000101010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--554
WHEN "0000001000101011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--555
WHEN "0000001000101100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--556
WHEN "0000001000101101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--557
WHEN "0000001000101110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--558
WHEN "0000001000101111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--559
WHEN "0000001000110000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--560
WHEN "0000001000110001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--561
WHEN "0000001000110010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--562
WHEN "0000001000110011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--563
WHEN "0000001000110100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--564
WHEN "0000001000110101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--565
WHEN "0000001000110110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--566
WHEN "0000001000110111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--567
WHEN "0000001000111000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--568
WHEN "0000001000111001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--569
WHEN "0000001000111010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--570
WHEN "0000001000111011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--571
WHEN "0000001000111100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--572
WHEN "0000001000111101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--573
WHEN "0000001000111110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--574
WHEN "0000001000111111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--575
WHEN "0000001001000000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--576
WHEN "0000001001000001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--577
WHEN "0000001001000010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--578
WHEN "0000001001000011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--579
WHEN "0000001001000100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--580
WHEN "0000001001000101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--581
WHEN "0000001001000110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--582
WHEN "0000001001000111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--583
WHEN "0000001001001000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--584
WHEN "0000001001001001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--585
WHEN "0000001001001010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--586
WHEN "0000001001001011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--587
WHEN "0000001001001100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--588
WHEN "0000001001001101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--589
WHEN "0000001001001110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--590
WHEN "0000001001001111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--591
WHEN "0000001001010000" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--592
WHEN "0000001001010001" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--593
WHEN "0000001001010010" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--594
WHEN "0000001001010011" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--595
WHEN "0000001001010100" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--596
WHEN "0000001001010101" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--597
WHEN "0000001001010110" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--598
WHEN "0000001001010111" => HEX3_D <= "1000000"; HEX2_D <= "0010010"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--599
WHEN "0000001001011000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--600
WHEN "0000001001011001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--601
WHEN "0000001001011010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--602
WHEN "0000001001011011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--603
WHEN "0000001001011100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--604
WHEN "0000001001011101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--605
WHEN "0000001001011110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--606
WHEN "0000001001011111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--607
WHEN "0000001001100000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--608
WHEN "0000001001100001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--609
WHEN "0000001001100010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--610
WHEN "0000001001100011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--611
WHEN "0000001001100100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--612
WHEN "0000001001100101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--613
WHEN "0000001001100110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--614
WHEN "0000001001100111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--615
WHEN "0000001001101000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--616
WHEN "0000001001101001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--617
WHEN "0000001001101010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--618
WHEN "0000001001101011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--619
WHEN "0000001001101100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--620
WHEN "0000001001101101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--621
WHEN "0000001001101110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--622
WHEN "0000001001101111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--623
WHEN "0000001001110000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--624
WHEN "0000001001110001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--625
WHEN "0000001001110010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--626
WHEN "0000001001110011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--627
WHEN "0000001001110100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--628
WHEN "0000001001110101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--629
WHEN "0000001001110110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--630
WHEN "0000001001110111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--631
WHEN "0000001001111000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--632
WHEN "0000001001111001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--633
WHEN "0000001001111010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--634
WHEN "0000001001111011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--635
WHEN "0000001001111100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--636
WHEN "0000001001111101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--637
WHEN "0000001001111110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--638
WHEN "0000001001111111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--639
WHEN "0000001010000000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--640
WHEN "0000001010000001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--641
WHEN "0000001010000010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--642
WHEN "0000001010000011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--643
WHEN "0000001010000100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--644
WHEN "0000001010000101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--645
WHEN "0000001010000110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--646
WHEN "0000001010000111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--647
WHEN "0000001010001000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--648
WHEN "0000001010001001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--649
WHEN "0000001010001010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--650
WHEN "0000001010001011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--651
WHEN "0000001010001100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--652
WHEN "0000001010001101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--653
WHEN "0000001010001110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--654
WHEN "0000001010001111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--655
WHEN "0000001010010000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--656
WHEN "0000001010010001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--657
WHEN "0000001010010010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--658
WHEN "0000001010010011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--659
WHEN "0000001010010100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--660
WHEN "0000001010010101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--661
WHEN "0000001010010110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--662
WHEN "0000001010010111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--663
WHEN "0000001010011000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--664
WHEN "0000001010011001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--665
WHEN "0000001010011010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--666
WHEN "0000001010011011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--667
WHEN "0000001010011100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--668
WHEN "0000001010011101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--669
WHEN "0000001010011110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--670
WHEN "0000001010011111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--671
WHEN "0000001010100000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--672
WHEN "0000001010100001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--673
WHEN "0000001010100010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--674
WHEN "0000001010100011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--675
WHEN "0000001010100100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--676
WHEN "0000001010100101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--677
WHEN "0000001010100110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--678
WHEN "0000001010100111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--679
WHEN "0000001010101000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--680
WHEN "0000001010101001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--681
WHEN "0000001010101010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--682
WHEN "0000001010101011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--683
WHEN "0000001010101100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--684
WHEN "0000001010101101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--685
WHEN "0000001010101110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--686
WHEN "0000001010101111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--687
WHEN "0000001010110000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--688
WHEN "0000001010110001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--689
WHEN "0000001010110010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--690
WHEN "0000001010110011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--691
WHEN "0000001010110100" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--692
WHEN "0000001010110101" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--693
WHEN "0000001010110110" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--694
WHEN "0000001010110111" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--695
WHEN "0000001010111000" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--696
WHEN "0000001010111001" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--697
WHEN "0000001010111010" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--698
WHEN "0000001010111011" => HEX3_D <= "1000000"; HEX2_D <= "0000010"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--699
WHEN "0000001010111100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--700
WHEN "0000001010111101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--701
WHEN "0000001010111110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--702
WHEN "0000001010111111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--703
WHEN "0000001011000000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--704
WHEN "0000001011000001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--705
WHEN "0000001011000010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--706
WHEN "0000001011000011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--707
WHEN "0000001011000100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--708
WHEN "0000001011000101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--709
WHEN "0000001011000110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--710
WHEN "0000001011000111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--711
WHEN "0000001011001000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--712
WHEN "0000001011001001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--713
WHEN "0000001011001010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--714
WHEN "0000001011001011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--715
WHEN "0000001011001100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--716
WHEN "0000001011001101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--717
WHEN "0000001011001110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--718
WHEN "0000001011001111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--719
WHEN "0000001011010000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--720
WHEN "0000001011010001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--721
WHEN "0000001011010010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--722
WHEN "0000001011010011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--723
WHEN "0000001011010100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--724
WHEN "0000001011010101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--725
WHEN "0000001011010110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--726
WHEN "0000001011010111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--727
WHEN "0000001011011000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--728
WHEN "0000001011011001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--729
WHEN "0000001011011010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--730
WHEN "0000001011011011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--731
WHEN "0000001011011100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--732
WHEN "0000001011011101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--733
WHEN "0000001011011110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--734
WHEN "0000001011011111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--735
WHEN "0000001011100000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--736
WHEN "0000001011100001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--737
WHEN "0000001011100010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--738
WHEN "0000001011100011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--739
WHEN "0000001011100100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--740
WHEN "0000001011100101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--741
WHEN "0000001011100110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--742
WHEN "0000001011100111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--743
WHEN "0000001011101000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--744
WHEN "0000001011101001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--745
WHEN "0000001011101010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--746
WHEN "0000001011101011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--747
WHEN "0000001011101100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--748
WHEN "0000001011101101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--749
WHEN "0000001011101110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--750
WHEN "0000001011101111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--751
WHEN "0000001011110000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--752
WHEN "0000001011110001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--753
WHEN "0000001011110010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--754
WHEN "0000001011110011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--755
WHEN "0000001011110100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--756
WHEN "0000001011110101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--757
WHEN "0000001011110110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--758
WHEN "0000001011110111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--759
WHEN "0000001011111000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--760
WHEN "0000001011111001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--761
WHEN "0000001011111010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--762
WHEN "0000001011111011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--763
WHEN "0000001011111100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--764
WHEN "0000001011111101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--765
WHEN "0000001011111110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--766
WHEN "0000001011111111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--767
WHEN "0000001100000000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--768
WHEN "0000001100000001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--769
WHEN "0000001100000010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--770
WHEN "0000001100000011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--771
WHEN "0000001100000100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--772
WHEN "0000001100000101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--773
WHEN "0000001100000110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--774
WHEN "0000001100000111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--775
WHEN "0000001100001000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--776
WHEN "0000001100001001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--777
WHEN "0000001100001010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--778
WHEN "0000001100001011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--779
WHEN "0000001100001100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--780
WHEN "0000001100001101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--781
WHEN "0000001100001110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--782
WHEN "0000001100001111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--783
WHEN "0000001100010000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--784
WHEN "0000001100010001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--785
WHEN "0000001100010010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--786
WHEN "0000001100010011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--787
WHEN "0000001100010100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--788
WHEN "0000001100010101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--789
WHEN "0000001100010110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--790
WHEN "0000001100010111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--791
WHEN "0000001100011000" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--792
WHEN "0000001100011001" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--793
WHEN "0000001100011010" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--794
WHEN "0000001100011011" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--795
WHEN "0000001100011100" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--796
WHEN "0000001100011101" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--797
WHEN "0000001100011110" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--798
WHEN "0000001100011111" => HEX3_D <= "1000000"; HEX2_D <= "1111000"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--799
WHEN "0000001100100000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--800
WHEN "0000001100100001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--801
WHEN "0000001100100010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--802
WHEN "0000001100100011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--803
WHEN "0000001100100100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--804
WHEN "0000001100100101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--805
WHEN "0000001100100110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--806
WHEN "0000001100100111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--807
WHEN "0000001100101000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--808
WHEN "0000001100101001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--809
WHEN "0000001100101010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--810
WHEN "0000001100101011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--811
WHEN "0000001100101100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--812
WHEN "0000001100101101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--813
WHEN "0000001100101110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--814
WHEN "0000001100101111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--815
WHEN "0000001100110000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--816
WHEN "0000001100110001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--817
WHEN "0000001100110010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--818
WHEN "0000001100110011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--819
WHEN "0000001100110100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--820
WHEN "0000001100110101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--821
WHEN "0000001100110110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--822
WHEN "0000001100110111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--823
WHEN "0000001100111000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--824
WHEN "0000001100111001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--825
WHEN "0000001100111010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--826
WHEN "0000001100111011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--827
WHEN "0000001100111100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--828
WHEN "0000001100111101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--829
WHEN "0000001100111110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--830
WHEN "0000001100111111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--831
WHEN "0000001101000000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--832
WHEN "0000001101000001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--833
WHEN "0000001101000010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--834
WHEN "0000001101000011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--835
WHEN "0000001101000100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--836
WHEN "0000001101000101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--837
WHEN "0000001101000110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--838
WHEN "0000001101000111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--839
WHEN "0000001101001000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--840
WHEN "0000001101001001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--841
WHEN "0000001101001010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--842
WHEN "0000001101001011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--843
WHEN "0000001101001100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--844
WHEN "0000001101001101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--845
WHEN "0000001101001110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--846
WHEN "0000001101001111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--847
WHEN "0000001101010000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--848
WHEN "0000001101010001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--849
WHEN "0000001101010010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--850
WHEN "0000001101010011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--851
WHEN "0000001101010100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--852
WHEN "0000001101010101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--853
WHEN "0000001101010110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--854
WHEN "0000001101010111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--855
WHEN "0000001101011000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--856
WHEN "0000001101011001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--857
WHEN "0000001101011010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--858
WHEN "0000001101011011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--859
WHEN "0000001101011100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--860
WHEN "0000001101011101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--861
WHEN "0000001101011110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--862
WHEN "0000001101011111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--863
WHEN "0000001101100000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--864
WHEN "0000001101100001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--865
WHEN "0000001101100010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--866
WHEN "0000001101100011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--867
WHEN "0000001101100100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--868
WHEN "0000001101100101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--869
WHEN "0000001101100110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--870
WHEN "0000001101100111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--871
WHEN "0000001101101000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--872
WHEN "0000001101101001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--873
WHEN "0000001101101010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--874
WHEN "0000001101101011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--875
WHEN "0000001101101100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--876
WHEN "0000001101101101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--877
WHEN "0000001101101110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--878
WHEN "0000001101101111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--879
WHEN "0000001101110000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--880
WHEN "0000001101110001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--881
WHEN "0000001101110010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--882
WHEN "0000001101110011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--883
WHEN "0000001101110100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--884
WHEN "0000001101110101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--885
WHEN "0000001101110110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--886
WHEN "0000001101110111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--887
WHEN "0000001101111000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--888
WHEN "0000001101111001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--889
WHEN "0000001101111010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--890
WHEN "0000001101111011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--891
WHEN "0000001101111100" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--892
WHEN "0000001101111101" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--893
WHEN "0000001101111110" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--894
WHEN "0000001101111111" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--895
WHEN "0000001110000000" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--896
WHEN "0000001110000001" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--897
WHEN "0000001110000010" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--898
WHEN "0000001110000011" => HEX3_D <= "1000000"; HEX2_D <= "0000000"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--899
WHEN "0000001110000100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--900
WHEN "0000001110000101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--901
WHEN "0000001110000110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--902
WHEN "0000001110000111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--903
WHEN "0000001110001000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--904
WHEN "0000001110001001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--905
WHEN "0000001110001010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--906
WHEN "0000001110001011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--907
WHEN "0000001110001100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--908
WHEN "0000001110001101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--909
WHEN "0000001110001110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--910
WHEN "0000001110001111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--911
WHEN "0000001110010000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--912
WHEN "0000001110010001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--913
WHEN "0000001110010010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--914
WHEN "0000001110010011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--915
WHEN "0000001110010100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--916
WHEN "0000001110010101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--917
WHEN "0000001110010110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--918
WHEN "0000001110010111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--919
WHEN "0000001110011000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--920
WHEN "0000001110011001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--921
WHEN "0000001110011010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--922
WHEN "0000001110011011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--923
WHEN "0000001110011100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0011001";--924
WHEN "0000001110011101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0010010";--925
WHEN "0000001110011110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0000010";--926
WHEN "0000001110011111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "1111000";--927
WHEN "0000001110100000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0000000";--928
WHEN "0000001110100001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0100100"; HEX0_D <= "0010000";--929
WHEN "0000001110100010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "1000000";--930
WHEN "0000001110100011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "1111001";--931
WHEN "0000001110100100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0100100";--932
WHEN "0000001110100101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0110000";--933
WHEN "0000001110100110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0011001";--934
WHEN "0000001110100111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0010010";--935
WHEN "0000001110101000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0000010";--936
WHEN "0000001110101001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "1111000";--937
WHEN "0000001110101010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0000000";--938
WHEN "0000001110101011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0110000"; HEX0_D <= "0010000";--939
WHEN "0000001110101100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "1000000";--940
WHEN "0000001110101101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "1111001";--941
WHEN "0000001110101110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0100100";--942
WHEN "0000001110101111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0110000";--943
WHEN "0000001110110000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0011001";--944
WHEN "0000001110110001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0010010";--945
WHEN "0000001110110010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0000010";--946
WHEN "0000001110110011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "1111000";--947
WHEN "0000001110110100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0000000";--948
WHEN "0000001110110101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0011001"; HEX0_D <= "0010000";--949
WHEN "0000001110110110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "1000000";--950
WHEN "0000001110110111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "1111001";--951
WHEN "0000001110111000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0100100";--952
WHEN "0000001110111001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0110000";--953
WHEN "0000001110111010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0011001";--954
WHEN "0000001110111011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0010010";--955
WHEN "0000001110111100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0000010";--956
WHEN "0000001110111101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "1111000";--957
WHEN "0000001110111110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0000000";--958
WHEN "0000001110111111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010010"; HEX0_D <= "0010000";--959
WHEN "0000001111000000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "1000000";--960
WHEN "0000001111000001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "1111001";--961
WHEN "0000001111000010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0100100";--962
WHEN "0000001111000011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0110000";--963
WHEN "0000001111000100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0011001";--964
WHEN "0000001111000101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0010010";--965
WHEN "0000001111000110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0000010";--966
WHEN "0000001111000111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "1111000";--967
WHEN "0000001111001000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0000000";--968
WHEN "0000001111001001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000010"; HEX0_D <= "0010000";--969
WHEN "0000001111001010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "1000000";--970
WHEN "0000001111001011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "1111001";--971
WHEN "0000001111001100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0100100";--972
WHEN "0000001111001101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0110000";--973
WHEN "0000001111001110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0011001";--974
WHEN "0000001111001111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0010010";--975
WHEN "0000001111010000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0000010";--976
WHEN "0000001111010001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "1111000";--977
WHEN "0000001111010010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0000000";--978
WHEN "0000001111010011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "1111000"; HEX0_D <= "0010000";--979
WHEN "0000001111010100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "1000000";--980
WHEN "0000001111010101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "1111001";--981
WHEN "0000001111010110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0100100";--982
WHEN "0000001111010111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0110000";--983
WHEN "0000001111011000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0011001";--984
WHEN "0000001111011001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0010010";--985
WHEN "0000001111011010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0000010";--986
WHEN "0000001111011011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "1111000";--987
WHEN "0000001111011100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0000000";--988
WHEN "0000001111011101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0000000"; HEX0_D <= "0010000";--989
WHEN "0000001111011110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "1000000";--990
WHEN "0000001111011111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "1111001";--991
WHEN "0000001111100000" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0100100";--992
WHEN "0000001111100001" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0110000";--993
WHEN "0000001111100010" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0011001";--994
WHEN "0000001111100011" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0010010";--995
WHEN "0000001111100100" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0000010";--996
WHEN "0000001111100101" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "1111000";--997
WHEN "0000001111100110" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0000000";--998
WHEN "0000001111100111" => HEX3_D <= "1000000"; HEX2_D <= "0010000"; HEX1_D <= "0010000"; HEX0_D <= "0010000";--999
WHEN "0000001111101000" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1000000";--1000
WHEN "0000001111101001" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1111001";--1001
WHEN "0000001111101010" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0100100";--1002
WHEN "0000001111101011" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0110000";--1003
WHEN "0000001111101100" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0011001";--1004
WHEN "0000001111101101" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0010010";--1005
WHEN "0000001111101110" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0000010";--1006
WHEN "0000001111101111" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "1111000";--1007
WHEN "0000001111110000" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0000000";--1008
WHEN "0000001111110001" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1000000"; HEX0_D <= "0010000";--1009
WHEN "0000001111110010" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1000000";--1010
WHEN "0000001111110011" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1111001";--1011
WHEN "0000001111110100" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0100100";--1012
WHEN "0000001111110101" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0110000";--1013
WHEN "0000001111110110" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0011001";--1014
WHEN "0000001111110111" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0010010";--1015
WHEN "0000001111111000" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0000010";--1016
WHEN "0000001111111001" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "1111000";--1017
WHEN "0000001111111010" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0000000";--1018
WHEN "0000001111111011" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "1111001"; HEX0_D <= "0010000";--1019
WHEN "0000001111111100" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "1000000";--1020
WHEN "0000001111111101" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "1111001";--1021
WHEN "0000001111111110" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0100100";--1022
WHEN "0000001111111111" => HEX3_D <= "1111001"; HEX2_D <= "1000000"; HEX1_D <= "0100100"; HEX0_D <= "0110000";--1023

WHEN OTHERS     => HEX3_D <= "0000110"; HEX2_D <= "0101011"; HEX1_D <= "0101011"; HEX0_D <= "0100011";
END CASE;
END IF;
END PROCESS;
END architecture;

